
module ByteSub_ShiftRow
(
  ap_clk,
  ap_rst,
  ap_start,
  ap_done,
  ap_idle,
  ap_ready,
  statemt_address0,
  statemt_ce0,
  statemt_we0,
  statemt_d0,
  statemt_q0,
  statemt_address1,
  statemt_ce1,
  statemt_we1,
  statemt_d1,
  statemt_q1,
  working_key
);

  parameter ap_ST_fsm_state1 = 16'd1;
  parameter ap_ST_fsm_state2 = 16'd2;
  parameter ap_ST_fsm_state3 = 16'd4;
  parameter ap_ST_fsm_state4 = 16'd8;
  parameter ap_ST_fsm_state5 = 16'd16;
  parameter ap_ST_fsm_state6 = 16'd32;
  parameter ap_ST_fsm_state7 = 16'd64;
  parameter ap_ST_fsm_state8 = 16'd128;
  parameter ap_ST_fsm_state9 = 16'd256;
  parameter ap_ST_fsm_state10 = 16'd512;
  parameter ap_ST_fsm_state11 = 16'd1024;
  parameter ap_ST_fsm_state12 = 16'd2048;
  parameter ap_ST_fsm_state13 = 16'd4096;
  parameter ap_ST_fsm_state14 = 16'd8192;
  parameter ap_ST_fsm_state15 = 16'd16384;
  parameter ap_ST_fsm_state16 = 16'd32768;
  input ap_clk;
  input ap_rst;
  input ap_start;
  output ap_done;
  output ap_idle;
  output ap_ready;
  output [4:0] statemt_address0;
  output statemt_ce0;
  output statemt_we0;
  output [31:0] statemt_d0;
  input [31:0] statemt_q0;
  output [4:0] statemt_address1;
  output statemt_ce1;
  output statemt_we1;
  output [31:0] statemt_d1;
  input [31:0] statemt_q1;
  reg ap_done;
  reg ap_idle;
  reg ap_ready;
  reg [4:0] statemt_address0;
  reg statemt_ce0;
  reg statemt_we0;
  reg [31:0] statemt_d0;
  reg [4:0] statemt_address1;
  reg statemt_ce1;
  reg statemt_we1;
  reg [31:0] statemt_d1;
  reg [15:0] ap_CS_fsm;
  wire ap_CS_fsm_state1;
  reg [7:0] Sbox_address0;
  reg Sbox_ce0;
  wire [7:0] Sbox_q0;
  reg [7:0] Sbox_address1;
  reg Sbox_ce1;
  wire [7:0] Sbox_q1;
  reg [7:0] reg_326;
  wire ap_CS_fsm_state3;
  wire ap_CS_fsm_state10;
  reg [7:0] reg_330;
  wire ap_CS_fsm_state9;
  reg [7:0] reg_335;
  wire ap_CS_fsm_state4;
  reg [7:0] reg_340;
  wire [4:0] statemt_addr_9_reg_496;
  wire [4:0] statemt_addr_10_reg_501;
  wire ap_CS_fsm_state2;
  wire [4:0] statemt_addr_11_reg_516;
  wire [4:0] statemt_addr_12_reg_521;
  wire [4:0] statemt_addr_13_reg_536;
  wire [4:0] statemt_addr_14_reg_541;
  wire [4:0] statemt_addr_15_reg_556;
  wire [4:0] statemt_addr_16_reg_561;
  reg [7:0] temp_1_reg_566;
  wire ap_CS_fsm_state5;
  reg [7:0] Sbox_load_4_reg_571;
  wire [4:0] statemt_addr_17_reg_586;
  wire [4:0] statemt_addr_18_reg_591;
  reg [7:0] temp_2_reg_596;
  wire ap_CS_fsm_state6;
  reg [7:0] Sbox_load_6_reg_601;
  wire [4:0] statemt_addr_19_reg_616;
  wire [4:0] statemt_addr_20_reg_621;
  wire [4:0] statemt_addr_reg_626;
  wire ap_CS_fsm_state7;
  reg [7:0] temp_3_reg_631;
  reg [7:0] Sbox_load_8_reg_636;
  wire [4:0] statemt_addr_21_reg_651;
  reg [7:0] Sbox_load_9_reg_656;
  wire ap_CS_fsm_state8;
  reg [7:0] Sbox_load_10_reg_661;
  wire [4:0] statemt_addr_22_reg_676;
  wire [4:0] statemt_addr_23_reg_681;
  wire signed [63:0] tmp_fu_344_p1;
  wire signed [63:0] tmp_s_fu_349_p1;
  wire signed [63:0] tmp_54_fu_354_p1;
  wire signed [63:0] tmp_55_fu_359_p1;
  wire signed [63:0] tmp_56_fu_364_p1;
  wire signed [63:0] tmp_57_fu_369_p1;
  wire signed [63:0] tmp_58_fu_374_p1;
  wire signed [63:0] tmp_59_fu_379_p1;
  wire signed [63:0] tmp_60_fu_384_p1;
  wire signed [63:0] tmp_61_fu_389_p1;
  wire signed [63:0] tmp_62_fu_394_p1;
  wire signed [63:0] tmp_63_fu_399_p1;
  wire signed [63:0] tmp_64_fu_404_p1;
  wire signed [63:0] tmp_65_fu_409_p1;
  wire signed [63:0] tmp_66_fu_424_p1;
  wire signed [63:0] tmp_67_fu_429_p1;
  wire [31:0] Sbox_load_cast_fu_414_p1;
  wire [31:0] Sbox_load_1_cast_fu_419_p1;
  wire [31:0] Sbox_load_2_cast_fu_439_p1;
  wire [31:0] temp_cast_fu_434_p1;
  wire ap_CS_fsm_state11;
  wire [31:0] Sbox_load_4_cast_fu_448_p1;
  wire [31:0] temp_1_cast_fu_444_p1;
  wire ap_CS_fsm_state12;
  wire [31:0] Sbox_load_6_cast_fu_456_p1;
  wire [31:0] temp_2_cast_fu_452_p1;
  wire ap_CS_fsm_state13;
  wire [31:0] Sbox_load_8_cast_fu_460_p1;
  wire [31:0] Sbox_load_9_cast_fu_464_p1;
  wire ap_CS_fsm_state14;
  wire [31:0] Sbox_load_10_cast_fu_472_p1;
  wire [31:0] temp_3_cast_fu_468_p1;
  wire ap_CS_fsm_state15;
  wire [31:0] Sbox_load_11_cast_fu_476_p1;
  wire [31:0] Sbox_load_12_cast_fu_481_p1;
  wire ap_CS_fsm_state16;
  wire [31:0] Sbox_load_13_cast_fu_486_p1;
  wire [31:0] Sbox_load_14_cast_fu_491_p1;
  wire signed [31:0] tmp_fu_344_p0;
  wire signed [31:0] tmp_s_fu_349_p0;
  wire signed [31:0] tmp_54_fu_354_p0;
  wire signed [31:0] tmp_55_fu_359_p0;
  wire signed [31:0] tmp_56_fu_364_p0;
  wire signed [31:0] tmp_57_fu_369_p0;
  wire signed [31:0] tmp_58_fu_374_p0;
  wire signed [31:0] tmp_59_fu_379_p0;
  wire signed [31:0] tmp_60_fu_384_p0;
  wire signed [31:0] tmp_61_fu_389_p0;
  wire signed [31:0] tmp_62_fu_394_p0;
  wire signed [31:0] tmp_63_fu_399_p0;
  wire signed [31:0] tmp_64_fu_404_p0;
  wire signed [31:0] tmp_65_fu_409_p0;
  wire signed [31:0] tmp_66_fu_424_p0;
  wire signed [31:0] tmp_67_fu_429_p0;
  reg [15:0] ap_NS_fsm;
  input [127:0] working_key;

  initial begin
    #0 ap_CS_fsm = 16'd1;
  end


  ByteSub_ShiftRow_bkb
  #(
    .DataWidth(8),
    .AddressRange(256),
    .AddressWidth(8)
  )
  Sbox_U
  (
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(Sbox_address0),
    .ce0(Sbox_ce0),
    .q0(Sbox_q0),
    .address1(Sbox_address1),
    .ce1(Sbox_ce1),
    .q1(Sbox_q1)
  );


  always @(posedge ap_clk) begin
    if(ap_rst == 1'b1) begin
      ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
      ap_CS_fsm <= ap_NS_fsm;
    end
  end


  always @(posedge ap_clk) begin
    if(1'b1 == ap_CS_fsm_state9) begin
      reg_330 <= Sbox_q0;
    end else if(1'b1 == ap_CS_fsm_state3) begin
      reg_330 <= Sbox_q1;
    end 
  end


  always @(posedge ap_clk) begin
    if(1'b1 == ap_CS_fsm_state9) begin
      reg_335 <= Sbox_q1;
    end else if(1'b1 == ap_CS_fsm_state4) begin
      reg_335 <= Sbox_q0;
    end 
  end


  always @(posedge ap_clk) begin
    if(1'b1 == ap_CS_fsm_state8) begin
      Sbox_load_10_reg_661 <= Sbox_q1;
      Sbox_load_9_reg_656 <= Sbox_q0;
    end 
  end


  always @(posedge ap_clk) begin
    if(1'b1 == ap_CS_fsm_state5) begin
      Sbox_load_4_reg_571 <= Sbox_q1;
      temp_1_reg_566 <= Sbox_q0;
    end 
  end


  always @(posedge ap_clk) begin
    if(1'b1 == ap_CS_fsm_state6) begin
      Sbox_load_6_reg_601 <= Sbox_q1;
      temp_2_reg_596 <= Sbox_q0;
    end 
  end


  always @(posedge ap_clk) begin
    if(1'b1 == ap_CS_fsm_state7) begin
      Sbox_load_8_reg_636 <= Sbox_q1;
      temp_3_reg_631 <= Sbox_q0;
    end 
  end


  always @(posedge ap_clk) begin
    if((1'b1 == ap_CS_fsm_state10) | (1'b1 == ap_CS_fsm_state3)) begin
      reg_326 <= Sbox_q0;
    end 
  end


  always @(posedge ap_clk) begin
    if((1'b1 == ap_CS_fsm_state4) | (1'b1 == ap_CS_fsm_state10)) begin
      reg_340 <= Sbox_q1;
    end 
  end


  always @(*) begin
    if(1'b1 == ap_CS_fsm_state9) begin
      Sbox_address0 = tmp_66_fu_424_p1;
    end else if(1'b1 == ap_CS_fsm_state8) begin
      Sbox_address0 = tmp_64_fu_404_p1;
    end else if(1'b1 == ap_CS_fsm_state7) begin
      Sbox_address0 = tmp_62_fu_394_p1;
    end else if(1'b1 == ap_CS_fsm_state6) begin
      Sbox_address0 = tmp_60_fu_384_p1;
    end else if(1'b1 == ap_CS_fsm_state5) begin
      Sbox_address0 = tmp_58_fu_374_p1;
    end else if(1'b1 == ap_CS_fsm_state4) begin
      Sbox_address0 = tmp_56_fu_364_p1;
    end else if(1'b1 == ap_CS_fsm_state3) begin
      Sbox_address0 = tmp_54_fu_354_p1;
    end else if(1'b1 == ap_CS_fsm_state2) begin
      Sbox_address0 = tmp_fu_344_p1;
    end else begin
      Sbox_address0 = 'bx;
    end
  end


  always @(*) begin
    if(1'b1 == ap_CS_fsm_state9) begin
      Sbox_address1 = tmp_67_fu_429_p1;
    end else if(1'b1 == ap_CS_fsm_state8) begin
      Sbox_address1 = tmp_65_fu_409_p1;
    end else if(1'b1 == ap_CS_fsm_state7) begin
      Sbox_address1 = tmp_63_fu_399_p1;
    end else if(1'b1 == ap_CS_fsm_state6) begin
      Sbox_address1 = tmp_61_fu_389_p1;
    end else if(1'b1 == ap_CS_fsm_state5) begin
      Sbox_address1 = tmp_59_fu_379_p1;
    end else if(1'b1 == ap_CS_fsm_state4) begin
      Sbox_address1 = tmp_57_fu_369_p1;
    end else if(1'b1 == ap_CS_fsm_state3) begin
      Sbox_address1 = tmp_55_fu_359_p1;
    end else if(1'b1 == ap_CS_fsm_state2) begin
      Sbox_address1 = tmp_s_fu_349_p1;
    end else begin
      Sbox_address1 = 'bx;
    end
  end


  always @(*) begin
    if((1'b1 == ap_CS_fsm_state2) | (1'b1 == ap_CS_fsm_state4) | (1'b1 == ap_CS_fsm_state9) | (1'b1 == ap_CS_fsm_state3) | (1'b1 == ap_CS_fsm_state8) | (1'b1 == ap_CS_fsm_state7) | (1'b1 == ap_CS_fsm_state6) | (1'b1 == ap_CS_fsm_state5)) begin
      Sbox_ce0 = 1'b1;
    end else begin
      Sbox_ce0 = 1'b0;
    end
  end


  always @(*) begin
    if((1'b1 == ap_CS_fsm_state2) | (1'b1 == ap_CS_fsm_state4) | (1'b1 == ap_CS_fsm_state9) | (1'b1 == ap_CS_fsm_state3) | (1'b1 == ap_CS_fsm_state8) | (1'b1 == ap_CS_fsm_state7) | (1'b1 == ap_CS_fsm_state6) | (1'b1 == ap_CS_fsm_state5)) begin
      Sbox_ce1 = 1'b1;
    end else begin
      Sbox_ce1 = 1'b0;
    end
  end


  always @(*) begin
    if((1'b1 == ap_CS_fsm_state16) | (ap_start == 1'b0) & (1'b1 == ap_CS_fsm_state1)) begin
      ap_done = 1'b1;
    end else begin
      ap_done = 1'b0;
    end
  end


  always @(*) begin
    if((ap_start == 1'b0) & (1'b1 == ap_CS_fsm_state1)) begin
      ap_idle = 1'b1;
    end else begin
      ap_idle = 1'b0;
    end
  end


  always @(*) begin
    if(1'b1 == ap_CS_fsm_state16) begin
      ap_ready = 1'b1;
    end else begin
      ap_ready = 1'b0;
    end
  end


  always @(*) begin
    if(1'b1 == ap_CS_fsm_state16) begin
      statemt_address0 = statemt_addr_22_reg_676;
    end else if(1'b1 == ap_CS_fsm_state15) begin
      statemt_address0 = statemt_addr_reg_626;
    end else if(1'b1 == ap_CS_fsm_state14) begin
      statemt_address0 = statemt_addr_19_reg_616;
    end else if(1'b1 == ap_CS_fsm_state13) begin
      statemt_address0 = statemt_addr_17_reg_586;
    end else if(1'b1 == ap_CS_fsm_state12) begin
      statemt_address0 = statemt_addr_15_reg_556;
    end else if(1'b1 == ap_CS_fsm_state11) begin
      statemt_address0 = statemt_addr_13_reg_536;
    end else if(1'b1 == ap_CS_fsm_state10) begin
      statemt_address0 = statemt_addr_11_reg_516;
    end else if(1'b1 == ap_CS_fsm_state9) begin
      statemt_address0 = statemt_addr_9_reg_496;
    end else if(1'b1 == ap_CS_fsm_state8) begin
      statemt_address0 = 64'd8;
    end else if(1'b1 == ap_CS_fsm_state7) begin
      statemt_address0 = 64'd0;
    end else if(1'b1 == ap_CS_fsm_state6) begin
      statemt_address0 = 64'd11;
    end else if(1'b1 == ap_CS_fsm_state5) begin
      statemt_address0 = 64'd3;
    end else if(1'b1 == ap_CS_fsm_state4) begin
      statemt_address0 = 64'd6;
    end else if(1'b1 == ap_CS_fsm_state3) begin
      statemt_address0 = 64'd2;
    end else if(1'b1 == ap_CS_fsm_state2) begin
      statemt_address0 = 64'd9;
    end else if(1'b1 == ap_CS_fsm_state1) begin
      statemt_address0 = 64'd1;
    end else begin
      statemt_address0 = 'bx;
    end
  end


  always @(*) begin
    if(1'b1 == ap_CS_fsm_state16) begin
      statemt_address1 = statemt_addr_23_reg_681;
    end else if(1'b1 == ap_CS_fsm_state15) begin
      statemt_address1 = statemt_addr_21_reg_651;
    end else if(1'b1 == ap_CS_fsm_state14) begin
      statemt_address1 = statemt_addr_20_reg_621;
    end else if(1'b1 == ap_CS_fsm_state13) begin
      statemt_address1 = statemt_addr_18_reg_591;
    end else if(1'b1 == ap_CS_fsm_state12) begin
      statemt_address1 = statemt_addr_16_reg_561;
    end else if(1'b1 == ap_CS_fsm_state11) begin
      statemt_address1 = statemt_addr_14_reg_541;
    end else if(1'b1 == ap_CS_fsm_state10) begin
      statemt_address1 = statemt_addr_12_reg_521;
    end else if(1'b1 == ap_CS_fsm_state9) begin
      statemt_address1 = statemt_addr_10_reg_501;
    end else if(1'b1 == ap_CS_fsm_state8) begin
      statemt_address1 = 64'd12;
    end else if(1'b1 == ap_CS_fsm_state7) begin
      statemt_address1 = 64'd4;
    end else if(1'b1 == ap_CS_fsm_state6) begin
      statemt_address1 = 64'd7;
    end else if(1'b1 == ap_CS_fsm_state5) begin
      statemt_address1 = 64'd15;
    end else if(1'b1 == ap_CS_fsm_state4) begin
      statemt_address1 = 64'd14;
    end else if(1'b1 == ap_CS_fsm_state3) begin
      statemt_address1 = 64'd10;
    end else if(1'b1 == ap_CS_fsm_state2) begin
      statemt_address1 = 64'd13;
    end else if(1'b1 == ap_CS_fsm_state1) begin
      statemt_address1 = 64'd5;
    end else begin
      statemt_address1 = 'bx;
    end
  end


  always @(*) begin
    if((1'b1 == ap_CS_fsm_state2) | (1'b1 == ap_CS_fsm_state4) | (1'b1 == ap_CS_fsm_state9) | (1'b1 == ap_CS_fsm_state10) | (1'b1 == ap_CS_fsm_state3) | (1'b1 == ap_CS_fsm_state16) | (1'b1 == ap_CS_fsm_state15) | (1'b1 == ap_CS_fsm_state14) | (1'b1 == ap_CS_fsm_state13) | (1'b1 == ap_CS_fsm_state12) | (1'b1 == ap_CS_fsm_state11) | (1'b1 == ap_CS_fsm_state8) | (1'b1 == ap_CS_fsm_state7) | (1'b1 == ap_CS_fsm_state6) | (1'b1 == ap_CS_fsm_state5) | (ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1)) begin
      statemt_ce0 = 1'b1;
    end else begin
      statemt_ce0 = 1'b0;
    end
  end


  always @(*) begin
    if((1'b1 == ap_CS_fsm_state2) | (1'b1 == ap_CS_fsm_state4) | (1'b1 == ap_CS_fsm_state9) | (1'b1 == ap_CS_fsm_state10) | (1'b1 == ap_CS_fsm_state3) | (1'b1 == ap_CS_fsm_state16) | (1'b1 == ap_CS_fsm_state15) | (1'b1 == ap_CS_fsm_state14) | (1'b1 == ap_CS_fsm_state13) | (1'b1 == ap_CS_fsm_state12) | (1'b1 == ap_CS_fsm_state11) | (1'b1 == ap_CS_fsm_state8) | (1'b1 == ap_CS_fsm_state7) | (1'b1 == ap_CS_fsm_state6) | (1'b1 == ap_CS_fsm_state5) | (ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1)) begin
      statemt_ce1 = 1'b1;
    end else begin
      statemt_ce1 = 1'b0;
    end
  end


  always @(*) begin
    if(1'b1 == ap_CS_fsm_state16) begin
      statemt_d0 = Sbox_load_13_cast_fu_486_p1;
    end else if(1'b1 == ap_CS_fsm_state15) begin
      statemt_d0 = Sbox_load_11_cast_fu_476_p1;
    end else if(1'b1 == ap_CS_fsm_state14) begin
      statemt_d0 = Sbox_load_10_cast_fu_472_p1;
    end else if(1'b1 == ap_CS_fsm_state13) begin
      statemt_d0 = Sbox_load_8_cast_fu_460_p1;
    end else if(1'b1 == ap_CS_fsm_state12) begin
      statemt_d0 = Sbox_load_6_cast_fu_456_p1;
    end else if(1'b1 == ap_CS_fsm_state11) begin
      statemt_d0 = Sbox_load_4_cast_fu_448_p1;
    end else if(1'b1 == ap_CS_fsm_state10) begin
      statemt_d0 = Sbox_load_2_cast_fu_439_p1;
    end else if(1'b1 == ap_CS_fsm_state9) begin
      statemt_d0 = Sbox_load_cast_fu_414_p1;
    end else begin
      statemt_d0 = 'bx;
    end
  end


  always @(*) begin
    if(1'b1 == ap_CS_fsm_state16) begin
      statemt_d1 = Sbox_load_14_cast_fu_491_p1;
    end else if(1'b1 == ap_CS_fsm_state15) begin
      statemt_d1 = Sbox_load_12_cast_fu_481_p1;
    end else if(1'b1 == ap_CS_fsm_state14) begin
      statemt_d1 = temp_3_cast_fu_468_p1;
    end else if(1'b1 == ap_CS_fsm_state13) begin
      statemt_d1 = Sbox_load_9_cast_fu_464_p1;
    end else if(1'b1 == ap_CS_fsm_state12) begin
      statemt_d1 = temp_2_cast_fu_452_p1;
    end else if(1'b1 == ap_CS_fsm_state11) begin
      statemt_d1 = temp_1_cast_fu_444_p1;
    end else if(1'b1 == ap_CS_fsm_state10) begin
      statemt_d1 = temp_cast_fu_434_p1;
    end else if(1'b1 == ap_CS_fsm_state9) begin
      statemt_d1 = Sbox_load_1_cast_fu_419_p1;
    end else begin
      statemt_d1 = 'bx;
    end
  end


  always @(*) begin
    if((1'b1 == ap_CS_fsm_state9) | (1'b1 == ap_CS_fsm_state10) | (1'b1 == ap_CS_fsm_state16) | (1'b1 == ap_CS_fsm_state15) | (1'b1 == ap_CS_fsm_state14) | (1'b1 == ap_CS_fsm_state13) | (1'b1 == ap_CS_fsm_state12) | (1'b1 == ap_CS_fsm_state11)) begin
      statemt_we0 = 1'b1;
    end else begin
      statemt_we0 = 1'b0;
    end
  end


  always @(*) begin
    if((1'b1 == ap_CS_fsm_state9) | (1'b1 == ap_CS_fsm_state10) | (1'b1 == ap_CS_fsm_state16) | (1'b1 == ap_CS_fsm_state15) | (1'b1 == ap_CS_fsm_state14) | (1'b1 == ap_CS_fsm_state13) | (1'b1 == ap_CS_fsm_state12) | (1'b1 == ap_CS_fsm_state11)) begin
      statemt_we1 = 1'b1;
    end else begin
      statemt_we1 = 1'b0;
    end
  end


  always @(*) begin
    case(ap_CS_fsm)
      ap_ST_fsm_state1: begin
        if((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1)) begin
          if(working_key[13] == 1'b1) begin
            ap_NS_fsm = ap_ST_fsm_state3;
          end else begin
            ap_NS_fsm = ap_ST_fsm_state2;
          end
        end else begin
          ap_NS_fsm = ap_ST_fsm_state1;
        end
      end
      ap_ST_fsm_state2: begin
        begin
          if(working_key[14] == 1'b1) begin
            ap_NS_fsm = ap_ST_fsm_state15;
          end else begin
            ap_NS_fsm = ap_ST_fsm_state3;
          end
        end
      end
      ap_ST_fsm_state3: begin
        begin
          if(working_key[15] == 1'b1) begin
            ap_NS_fsm = ap_ST_fsm_state5;
          end else begin
            ap_NS_fsm = ap_ST_fsm_state4;
          end
        end
      end
      ap_ST_fsm_state4: begin
        begin
          if(working_key[16] == 1'b1) begin
            ap_NS_fsm = ap_ST_fsm_state6;
          end else begin
            ap_NS_fsm = ap_ST_fsm_state5;
          end
        end
      end
      ap_ST_fsm_state5: begin
        begin
          if(working_key[17] == 1'b1) begin
            ap_NS_fsm = ap_ST_fsm_state15;
          end else begin
            ap_NS_fsm = ap_ST_fsm_state6;
          end
        end
      end
      ap_ST_fsm_state6: begin
        begin
          if(working_key[18] == 1'b1) begin
            ap_NS_fsm = ap_ST_fsm_state8;
          end else begin
            ap_NS_fsm = ap_ST_fsm_state7;
          end
        end
      end
      ap_ST_fsm_state7: begin
        begin
          if(working_key[19] == 1'b1) begin
            ap_NS_fsm = ap_ST_fsm_state9;
          end else begin
            ap_NS_fsm = ap_ST_fsm_state8;
          end
        end
      end
      ap_ST_fsm_state8: begin
        begin
          if(working_key[20] == 1'b1) begin
            ap_NS_fsm = ap_ST_fsm_state13;
          end else begin
            ap_NS_fsm = ap_ST_fsm_state9;
          end
        end
      end
      ap_ST_fsm_state9: begin
        begin
          if(working_key[21] == 1'b1) begin
            ap_NS_fsm = ap_ST_fsm_state14;
          end else begin
            ap_NS_fsm = ap_ST_fsm_state10;
          end
        end
      end
      ap_ST_fsm_state10: begin
        begin
          if(working_key[22] == 1'b1) begin
            ap_NS_fsm = ap_ST_fsm_state12;
          end else begin
            ap_NS_fsm = ap_ST_fsm_state11;
          end
        end
      end
      ap_ST_fsm_state11: begin
        begin
          if(working_key[23] == 1'b1) begin
            ap_NS_fsm = ap_ST_fsm_state15;
          end else begin
            ap_NS_fsm = ap_ST_fsm_state12;
          end
        end
      end
      ap_ST_fsm_state12: begin
        begin
          if(working_key[24] == 1'b1) begin
            ap_NS_fsm = ap_ST_fsm_state16;
          end else begin
            ap_NS_fsm = ap_ST_fsm_state13;
          end
        end
      end
      ap_ST_fsm_state13: begin
        ap_NS_fsm = ap_ST_fsm_state14;
      end
      ap_ST_fsm_state14: begin
        ap_NS_fsm = ap_ST_fsm_state15;
      end
      ap_ST_fsm_state15: begin
        ap_NS_fsm = ap_ST_fsm_state16;
      end
      ap_ST_fsm_state16: begin
        ap_NS_fsm = ap_ST_fsm_state1;
      end
      default: begin
        ap_NS_fsm = 'bx;
      end
    endcase
  end

  assign Sbox_load_10_cast_fu_472_p1 = Sbox_load_10_reg_661;
  assign Sbox_load_11_cast_fu_476_p1 = reg_330;
  assign Sbox_load_12_cast_fu_481_p1 = reg_335;
  assign Sbox_load_13_cast_fu_486_p1 = reg_326;
  assign Sbox_load_14_cast_fu_491_p1 = reg_340;
  assign Sbox_load_1_cast_fu_419_p1 = reg_335;
  assign Sbox_load_2_cast_fu_439_p1 = reg_340;
  assign Sbox_load_4_cast_fu_448_p1 = Sbox_load_4_reg_571;
  assign Sbox_load_6_cast_fu_456_p1 = Sbox_load_6_reg_601;
  assign Sbox_load_8_cast_fu_460_p1 = Sbox_load_8_reg_636;
  assign Sbox_load_9_cast_fu_464_p1 = Sbox_load_9_reg_656;
  assign Sbox_load_cast_fu_414_p1 = reg_330;
  assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];
  assign ap_CS_fsm_state10 = ap_CS_fsm[32'd9];
  assign ap_CS_fsm_state11 = ap_CS_fsm[32'd10];
  assign ap_CS_fsm_state12 = ap_CS_fsm[32'd11];
  assign ap_CS_fsm_state13 = ap_CS_fsm[32'd12];
  assign ap_CS_fsm_state14 = ap_CS_fsm[32'd13];
  assign ap_CS_fsm_state15 = ap_CS_fsm[32'd14];
  assign ap_CS_fsm_state16 = ap_CS_fsm[32'd15];
  assign ap_CS_fsm_state2 = ap_CS_fsm[32'd1];
  assign ap_CS_fsm_state3 = ap_CS_fsm[32'd2];
  assign ap_CS_fsm_state4 = ap_CS_fsm[32'd3];
  assign ap_CS_fsm_state5 = ap_CS_fsm[32'd4];
  assign ap_CS_fsm_state6 = ap_CS_fsm[32'd5];
  assign ap_CS_fsm_state7 = ap_CS_fsm[32'd6];
  assign ap_CS_fsm_state8 = ap_CS_fsm[32'd7];
  assign ap_CS_fsm_state9 = ap_CS_fsm[32'd8];
  assign statemt_addr_10_reg_501 = 64'd5;
  assign statemt_addr_11_reg_516 = 64'd9;
  assign statemt_addr_12_reg_521 = 64'd13;
  assign statemt_addr_13_reg_536 = 64'd2;
  assign statemt_addr_14_reg_541 = 64'd10;
  assign statemt_addr_15_reg_556 = 64'd6;
  assign statemt_addr_16_reg_561 = 64'd14;
  assign statemt_addr_17_reg_586 = 64'd3;
  assign statemt_addr_18_reg_591 = 64'd15;
  assign statemt_addr_19_reg_616 = 64'd11;
  assign statemt_addr_20_reg_621 = 64'd7;
  assign statemt_addr_21_reg_651 = 64'd4;
  assign statemt_addr_22_reg_676 = 64'd8;
  assign statemt_addr_23_reg_681 = 64'd12;
  assign statemt_addr_9_reg_496 = 64'd1;
  assign statemt_addr_reg_626 = 64'd0;
  assign temp_1_cast_fu_444_p1 = temp_1_reg_566;
  assign temp_2_cast_fu_452_p1 = temp_2_reg_596;
  assign temp_3_cast_fu_468_p1 = temp_3_reg_631;
  assign temp_cast_fu_434_p1 = reg_326;
  assign tmp_54_fu_354_p0 = statemt_q0;
  assign tmp_54_fu_354_p1 = tmp_54_fu_354_p0;
  assign tmp_55_fu_359_p0 = statemt_q1;
  assign tmp_55_fu_359_p1 = tmp_55_fu_359_p0;
  assign tmp_56_fu_364_p0 = statemt_q0;
  assign tmp_56_fu_364_p1 = tmp_56_fu_364_p0;
  assign tmp_57_fu_369_p0 = statemt_q1;
  assign tmp_57_fu_369_p1 = tmp_57_fu_369_p0;
  assign tmp_58_fu_374_p0 = statemt_q0;
  assign tmp_58_fu_374_p1 = tmp_58_fu_374_p0;
  assign tmp_59_fu_379_p0 = statemt_q1;
  assign tmp_59_fu_379_p1 = tmp_59_fu_379_p0;
  assign tmp_60_fu_384_p0 = statemt_q0;
  assign tmp_60_fu_384_p1 = tmp_60_fu_384_p0;
  assign tmp_61_fu_389_p0 = statemt_q1;
  assign tmp_61_fu_389_p1 = tmp_61_fu_389_p0;
  assign tmp_62_fu_394_p0 = statemt_q0;
  assign tmp_62_fu_394_p1 = tmp_62_fu_394_p0;
  assign tmp_63_fu_399_p0 = statemt_q1;
  assign tmp_63_fu_399_p1 = tmp_63_fu_399_p0;
  assign tmp_64_fu_404_p0 = statemt_q0;
  assign tmp_64_fu_404_p1 = tmp_64_fu_404_p0;
  assign tmp_65_fu_409_p0 = statemt_q1;
  assign tmp_65_fu_409_p1 = tmp_65_fu_409_p0;
  assign tmp_66_fu_424_p0 = statemt_q0;
  assign tmp_66_fu_424_p1 = tmp_66_fu_424_p0;
  assign tmp_67_fu_429_p0 = statemt_q1;
  assign tmp_67_fu_429_p1 = tmp_67_fu_429_p0;
  assign tmp_fu_344_p0 = statemt_q0;
  assign tmp_fu_344_p1 = tmp_fu_344_p0;
  assign tmp_s_fu_349_p0 = statemt_q1;
  assign tmp_s_fu_349_p1 = tmp_s_fu_349_p0;

endmodule

