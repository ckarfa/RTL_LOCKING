
module top_main
(
  ap_clk,
  ap_rst,
  ap_start,
  ap_done,
  ap_idle,
  ap_ready,
  ap_return,
  working_key
);

  parameter ap_ST_fsm_state1 = 6'd1;
  parameter ap_ST_fsm_state2 = 6'd2;
  parameter ap_ST_fsm_state3 = 6'd4;
  parameter ap_ST_fsm_state4 = 6'd8;
  parameter ap_ST_fsm_state5 = 6'd16;
  parameter ap_ST_fsm_state6 = 6'd32;
  input ap_clk;
  input ap_rst;
  input ap_start;
  output ap_done;
  output ap_idle;
  output ap_ready;
  output [31:0] ap_return;
  reg ap_done;
  reg ap_idle;
  reg ap_ready;
  reg [5:0] ap_CS_fsm;
  wire ap_CS_fsm_state1;
  wire [4:0] a_input_address0;
  reg a_input_ce0;
  wire [63:0] a_input_q0;
  wire [4:0] b_input_address0;
  reg b_input_ce0;
  wire [63:0] b_input_q0;
  wire [4:0] z_output_address0;
  reg z_output_ce0;
  wire [63:0] z_output_q0;
  wire [4:0] i_1_fu_128_p2;
  reg [4:0] i_1_reg_185;
  wire ap_CS_fsm_state2;
  wire [63:0] tmp_fu_134_p1;
  reg [63:0] tmp_reg_190;
  wire [0:0] exitcond_fu_122_p2;
  reg [63:0] x1_reg_205;
  wire ap_CS_fsm_state3;
  reg [63:0] x2_reg_210;
  wire [0:0] tmp_2_fu_144_p3;
  reg [0:0] tmp_2_reg_215;
  wire [0:0] tmp_itmp_fu_160_p2;
  reg [0:0] tmp_itmp_reg_220;
  wire [63:0] grp_subFloat64Sigs_fu_111_ap_return;
  wire ap_CS_fsm_state5;
  wire grp_subFloat64Sigs_fu_111_ap_ready;
  wire grp_subFloat64Sigs_fu_111_ap_done;
  reg ap_block_state5_on_subcall_done;
  wire [4:0] main_result_1_fu_176_p2;
  wire ap_CS_fsm_state6;
  wire grp_subFloat64Sigs_fu_111_ap_start;
  wire grp_subFloat64Sigs_fu_111_ap_idle;
  reg [4:0] i_reg_77;
  reg [4:0] main_result_reg_88;
  reg [63:0] result_reg_100;
  reg grp_subFloat64Sigs_fu_111_ap_start_reg;
  wire ap_CS_fsm_state4;
  wire [0:0] tmp_3_fu_152_p3;
  wire [0:0] tmp_1_fu_166_p2;
  wire [4:0] tmp_2_cast_fu_172_p1;
  reg [5:0] ap_NS_fsm;
  input [128:0] working_key;

  initial begin
    #0 ap_CS_fsm = 6'd1;
    #0 grp_subFloat64Sigs_fu_111_ap_start_reg = 1'b0;
  end


  top_main_a_input
  #(
    .DataWidth(64),
    .AddressRange(22),
    .AddressWidth(5)
  )
  a_input_U
  (
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(a_input_address0),
    .ce0(a_input_ce0),
    .q0(a_input_q0)
  );


  top_main_b_input
  #(
    .DataWidth(64),
    .AddressRange(22),
    .AddressWidth(5)
  )
  b_input_U
  (
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(b_input_address0),
    .ce0(b_input_ce0),
    .q0(b_input_q0)
  );


  top_main_z_output
  #(
    .DataWidth(64),
    .AddressRange(22),
    .AddressWidth(5)
  )
  z_output_U
  (
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(z_output_address0),
    .ce0(z_output_ce0),
    .q0(z_output_q0)
  );


  subFloat64Sigs
  grp_subFloat64Sigs_fu_111
  (
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(grp_subFloat64Sigs_fu_111_ap_start),
    .ap_done(grp_subFloat64Sigs_fu_111_ap_done),
    .ap_idle(grp_subFloat64Sigs_fu_111_ap_idle),
    .ap_ready(grp_subFloat64Sigs_fu_111_ap_ready),
    .a(x1_reg_205),
    .b(x2_reg_210),
    .zSign(tmp_2_reg_215),
    .ap_return(grp_subFloat64Sigs_fu_111_ap_return),
    .working_key(working_key)
  );


  always @(posedge ap_clk) begin
    if(ap_rst == 1'b1) begin
      ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
      ap_CS_fsm <= ap_NS_fsm;
    end
  end


  always @(posedge ap_clk) begin
    if(ap_rst == 1'b1) begin
      grp_subFloat64Sigs_fu_111_ap_start_reg <= 1'b0;
    end else begin
      if(1'b1 == ap_CS_fsm_state4) begin
        grp_subFloat64Sigs_fu_111_ap_start_reg <= 1'b1;
      end else if(grp_subFloat64Sigs_fu_111_ap_ready == 1'b1) begin
        grp_subFloat64Sigs_fu_111_ap_start_reg <= 1'b0;
      end 
    end
  end


  always @(posedge ap_clk) begin
    if(1'b1 == ap_CS_fsm_state6) begin
      if(working_key[0] == 1'b1) begin
        i_reg_77 <= a_input_q0;
      end else begin
        i_reg_77 <= i_1_reg_185;
      end
    end else if((1'b1 == ap_CS_fsm_state1) & (ap_start == 1'b1)) begin
      i_reg_77 <= 5'd0;
    end 
  end


  always @(posedge ap_clk) begin
    if(1'b1 == ap_CS_fsm_state6) begin
      if(working_key[1] == 1'b1) begin
        main_result_reg_88 <= main_result_1_fu_176_p2;
      end else begin
        main_result_reg_88 <= a_input_q0;
      end
    end else if((1'b1 == ap_CS_fsm_state1) & (ap_start == 1'b1)) begin
      main_result_reg_88 <= 5'd0;
    end 
  end


  always @(posedge ap_clk) begin
    if(1'b1 == ap_CS_fsm_state2) begin
      if(working_key[2] == 1'b1) begin
        i_1_reg_185 <= b_input_q0;
      end else begin
        i_1_reg_185 <= i_1_fu_128_p2;
      end
    end 
  end


  always @(posedge ap_clk) begin
    if((1'b0 == ap_block_state5_on_subcall_done) & (tmp_itmp_reg_220 == 1'd1) & (1'b1 == ap_CS_fsm_state5)) begin
      result_reg_100 <= grp_subFloat64Sigs_fu_111_ap_return;
    end 
  end


  always @(posedge ap_clk) begin
    if(1'b1 == ap_CS_fsm_state3) begin
      tmp_2_reg_215 <= a_input_q0[32'd63];
      tmp_itmp_reg_220 <= tmp_itmp_fu_160_p2;
      x1_reg_205 <= a_input_q0;
      x2_reg_210 <= b_input_q0;
    end 
  end


  always @(posedge ap_clk) begin
    if((exitcond_fu_122_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state2)) begin
      tmp_reg_190[4:0] <= tmp_fu_134_p1[4:0];
    end 
  end


  always @(*) begin
    if(1'b1 == ap_CS_fsm_state2) begin
      a_input_ce0 = 1'b1;
    end else begin
      a_input_ce0 = 1'b0;
    end
  end


  always @(*) begin
    if((exitcond_fu_122_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state2)) begin
      ap_done = 1'b1;
    end else begin
      ap_done = 1'b0;
    end
  end


  always @(*) begin
    if((ap_start == 1'b0) & (1'b1 == ap_CS_fsm_state1)) begin
      ap_idle = 1'b1;
    end else begin
      ap_idle = 1'b0;
    end
  end


  always @(*) begin
    if((exitcond_fu_122_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state2)) begin
      ap_ready = 1'b1;
    end else begin
      ap_ready = 1'b0;
    end
  end


  always @(*) begin
    if(1'b1 == ap_CS_fsm_state2) begin
      b_input_ce0 = 1'b1;
    end else begin
      b_input_ce0 = 1'b0;
    end
  end


  always @(*) begin
    if((1'b0 == ap_block_state5_on_subcall_done) & (1'b1 == ap_CS_fsm_state5)) begin
      z_output_ce0 = 1'b1;
    end else begin
      z_output_ce0 = 1'b0;
    end
  end


  always @(*) begin
    case(ap_CS_fsm)
      ap_ST_fsm_state1: begin
        if((1'b1 == ap_CS_fsm_state1) & (ap_start == 1'b1)) begin
          ap_NS_fsm = ap_ST_fsm_state2;
        end else begin
          ap_NS_fsm = ap_ST_fsm_state1;
        end
      end
      ap_ST_fsm_state2: begin
        if((exitcond_fu_122_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state2)) begin
          ap_NS_fsm = ap_ST_fsm_state1;
        end else begin
          ap_NS_fsm = ap_ST_fsm_state3;
        end
      end
      ap_ST_fsm_state3: begin
        if((tmp_itmp_fu_160_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state3)) begin
          ap_NS_fsm = ap_ST_fsm_state5;
        end else begin
          ap_NS_fsm = ap_ST_fsm_state4;
        end
      end
      ap_ST_fsm_state4: begin
        ap_NS_fsm = ap_ST_fsm_state5;
      end
      ap_ST_fsm_state5: begin
        if((1'b0 == ap_block_state5_on_subcall_done) & (1'b1 == ap_CS_fsm_state5)) begin
          ap_NS_fsm = ap_ST_fsm_state6;
        end else begin
          ap_NS_fsm = ap_ST_fsm_state5;
        end
      end
      ap_ST_fsm_state6: begin
        ap_NS_fsm = ap_ST_fsm_state2;
      end
      default: begin
        ap_NS_fsm = 'bx;
      end
    endcase
  end

  assign a_input_address0 = tmp_fu_134_p1;
  assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];
  assign ap_CS_fsm_state2 = ap_CS_fsm[32'd1];
  assign ap_CS_fsm_state3 = ap_CS_fsm[32'd2];
  assign ap_CS_fsm_state4 = ap_CS_fsm[32'd3];
  assign ap_CS_fsm_state5 = ap_CS_fsm[32'd4];
  assign ap_CS_fsm_state6 = ap_CS_fsm[32'd5];

  always @(*) begin
    ap_block_state5_on_subcall_done = (tmp_itmp_reg_220 == 1'd1) & (grp_subFloat64Sigs_fu_111_ap_done == 1'b0);
  end

  assign ap_return = main_result_reg_88;
  assign b_input_address0 = tmp_fu_134_p1;
  assign exitcond_fu_122_p2 = (i_reg_77 == 5'd22)? 1'b1 : 1'b0;
  assign grp_subFloat64Sigs_fu_111_ap_start = grp_subFloat64Sigs_fu_111_ap_start_reg;
  assign i_1_fu_128_p2 = i_reg_77 + 5'd1;
  assign main_result_1_fu_176_p2 = tmp_2_cast_fu_172_p1 + main_result_reg_88;
  assign tmp_1_fu_166_p2 = (result_reg_100 != z_output_q0)? 1'b1 : 1'b0;
  assign tmp_2_cast_fu_172_p1 = tmp_1_fu_166_p2;
  assign tmp_2_fu_144_p3 = a_input_q0[32'd63];
  assign tmp_3_fu_152_p3 = b_input_q0[32'd63];
  assign tmp_fu_134_p1 = i_reg_77;
  assign tmp_itmp_fu_160_p2 = tmp_3_fu_152_p3 ^ tmp_2_fu_144_p3;
  assign z_output_address0 = tmp_reg_190;

  always @(posedge ap_clk) begin
    tmp_reg_190[63:5] <= 59'b00000000000000000000000000000000000000000000000000000000000;
  end


endmodule

